`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 26.07.2025 18:45:59
// Design Name: 
// Module Name: fsm_lockout
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fsm_lockout;


    // Inputs
    reg clk;
    reg reset;
    reg [3:0] digit;
    reg enter;
    reg view_pass;
    reg set_pass;

    // Outputs
    wire green_led;
    wire red_led;
    wire alarm;
    wire [15:0] viewed_pass;
    wire [1:0] attempts_left;

    // DUT Instantiation
    fsm_password_lock dut (
        .clk(clk),
        .reset(reset),
        .digit(digit),
        .enter(enter),
        .view_pass(view_pass),
        .set_pass(set_pass),
        .green_led(green_led),
        .red_led(red_led),
        .alarm(alarm),
        .viewed_pass(viewed_pass),
        .attempts_left(attempts_left)
    );

    // Clock Generation
    always #5 clk = ~clk;

    // Task to input one digit
    task enter_digit(input [3:0] d);
    begin
        @(posedge clk);
        digit = d;
        enter = 1;
        @(posedge clk);
        enter = 0;
    end
    endtask

    // Task to enter 4-digit password
    task enter_password(input [3:0] d0, d1, d2, d3);
    begin
        enter_digit(d0);
        enter_digit(d1);
        enter_digit(d2);
        enter_digit(d3);
    end
    endtask

    initial begin
        // Init
        clk = 0;
        reset = 1;
        digit = 0;
        enter = 0;
        set_pass = 0;
        view_pass = 0;

        // Apply reset
        #10 reset = 0;

        // Attempt 1 - wrong password
        enter_password(9, 9, 9, 9);
        #40;

        // Attempt 2 - wrong password
        enter_password(8, 8, 8, 8);
        #40;

        // Attempt 3 - wrong password
        enter_password(7, 7, 7, 7);
        #60;

        // Check lockout condition
        $display("\n--- After 3 Wrong Attempts ---");
        $display("Alarm = %b | Red LED = %b | Green LED = %b | Attempts Left = %d",
                  alarm, red_led, green_led, attempts_left);

        // Try entering correct password after lockout
        enter_password(1, 2, 3, 4);  // default correct password
        #60;

        $display("\n--- After Trying Correct Password After Lockout ---");
        $display("Alarm = %b | Red LED = %b | Green LED = %b | Attempts Left = %d",
                  alarm, red_led, green_led, attempts_left);

        #20;
        $finish;
    end

    // Monitor internal state
    always @(posedge clk) begin
        $display("T=%0t | State=%0d | Digit=%h | Attempts=%d | Green=%b | Red=%b | Alarm=%b", 
                 $time, dut.curr_state, digit, attempts_left, green_led, red_led, alarm);
    end

endmodule


    

